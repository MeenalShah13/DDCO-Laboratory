module fa (input wire i0, i1, cin, output wire sum, cout); 
wire t0, t1, t2; 
xor3 _i0 (i0,i1,cin,sum);  
and2 _i1 (i0,i1,t0);   
and2 _i2 (i1,cin,t1); 
and2 _i3 (cin,i0,t2);  
or3 _i4 (t0,t1,t2,cout);
endmodule
