module p1(a,b,c,y);
input(a,b,c);
output(y);
wire(e,d);
and g1(e,a,b);
not g2(d,c);
or(y,e,d);
endmodule
